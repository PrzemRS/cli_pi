module licznik_gate(clk, nRst, led, ts_si, ts_so, scan_en);
  input  [0:0] ts_si;
  input  clk, nRst, scan_en;
  output [3:0] led;
  output [0:0] ts_so;

  wire clk_o, N2, N3, N4, n2, n6, n7, n8, n9, n10,
       ts_lockup_latchn_clkc0_intno3_, ts_pbuf_intsi37_;

  assign ts_so = ts_lockup_latchn_clkc0_intno3_;
  sffr \counter_reg[0] (
      .D(n2), .SI(ts_pbuf_intsi37_), .SE(scan_en), .CLK(clk_o), .R(n10), .Q(led[0]),
      .QB(n2)
  );
  sffr \counter_reg[1] (
      .D(N2), .SI(led[0]), .SE(scan_en), .CLK(clk_o), .R(n10), .Q(led[1]), .QB(n9)
  );
  sffr \counter_reg[2] (
      .D(N3), .SI(led[1]), .SE(scan_en), .CLK(clk_o), .R(n10), .Q(led[2]), .QB()
  );
  sffr \counter_reg[3] (
      .D(N4), .SI(led[2]), .SE(scan_en), .CLK(clk_o), .R(n10), .Q(led[3]), .QB(n8)
  );
  clock_divider2 clock_divider_inst(
      .clk_i(clk), .rst_i(nRst), .clk_o(clk_o)
  );
  inv01 U10(
      .A(nRst), .Y(n10)
  );
  xnor2 U11(
      .A0(n8), .A1(n6), .Y(N4)
  );
  nor02 U12(
      .A0(n7), .A1(led[2]), .Y(n6)
  );
  xnor2 U13(
      .A0(led[2]), .A1(n7), .Y(N3)
  );
  oai21 U14(
      .A0(n9), .A1(n2), .B0(n7), .Y(N2)
  );
  nand02 U15(
      .A0(n9), .A1(n2), .Y(n7)
  );
  nlatch ts_lockup_latchn_clkc0_intno3_i(
      .D(led[3]), .CLK(clk), .Q(ts_lockup_latchn_clkc0_intno3_)
  );
  buf02 tessent_persistent_cell_buf_intsi37_i(
      .A(ts_si), .Y(ts_pbuf_intsi37_)
  );
endmodule

/* Generated by Tessent Shell 2018.4-snapshot_2018.09.25_03.00 at Tue Sep 25 00:26:12 PDT 2018 */
module clock_divider_DW01_inc_0(A, SUM);
  input  [31:0] A;
  output [31:0] SUM;

  wire [31:2] carry;

  hadd1 \G1/G1_1(30)/U1_1 (
      .A(A[30]), .B(carry[30]), .S(SUM[30]), .CO(carry[31])
  );
  hadd1 \G1/G1_1(29)/U1_1 (
      .A(A[29]), .B(carry[29]), .S(SUM[29]), .CO(carry[30])
  );
  hadd1 \G1/G1_1(28)/U1_1 (
      .A(A[28]), .B(carry[28]), .S(SUM[28]), .CO(carry[29])
  );
  hadd1 \G1/G1_1(27)/U1_1 (
      .A(A[27]), .B(carry[27]), .S(SUM[27]), .CO(carry[28])
  );
  hadd1 \G1/G1_1(26)/U1_1 (
      .A(A[26]), .B(carry[26]), .S(SUM[26]), .CO(carry[27])
  );
  hadd1 \G1/G1_1(25)/U1_1 (
      .A(A[25]), .B(carry[25]), .S(SUM[25]), .CO(carry[26])
  );
  hadd1 \G1/G1_1(24)/U1_1 (
      .A(A[24]), .B(carry[24]), .S(SUM[24]), .CO(carry[25])
  );
  hadd1 \G1/G1_1(23)/U1_1 (
      .A(A[23]), .B(carry[23]), .S(SUM[23]), .CO(carry[24])
  );
  hadd1 \G1/G1_1(22)/U1_1 (
      .A(A[22]), .B(carry[22]), .S(SUM[22]), .CO(carry[23])
  );
  hadd1 \G1/G1_1(21)/U1_1 (
      .A(A[21]), .B(carry[21]), .S(SUM[21]), .CO(carry[22])
  );
  hadd1 \G1/G1_1(20)/U1_1 (
      .A(A[20]), .B(carry[20]), .S(SUM[20]), .CO(carry[21])
  );
  hadd1 \G1/G1_1(19)/U1_1 (
      .A(A[19]), .B(carry[19]), .S(SUM[19]), .CO(carry[20])
  );
  hadd1 \G1/G1_1(18)/U1_1 (
      .A(A[18]), .B(carry[18]), .S(SUM[18]), .CO(carry[19])
  );
  hadd1 \G1/G1_1(17)/U1_1 (
      .A(A[17]), .B(carry[17]), .S(SUM[17]), .CO(carry[18])
  );
  hadd1 \G1/G1_1(16)/U1_1 (
      .A(A[16]), .B(carry[16]), .S(SUM[16]), .CO(carry[17])
  );
  hadd1 \G1/G1_1(15)/U1_1 (
      .A(A[15]), .B(carry[15]), .S(SUM[15]), .CO(carry[16])
  );
  hadd1 \G1/G1_1(14)/U1_1 (
      .A(A[14]), .B(carry[14]), .S(SUM[14]), .CO(carry[15])
  );
  hadd1 \G1/G1_1(13)/U1_1 (
      .A(A[13]), .B(carry[13]), .S(SUM[13]), .CO(carry[14])
  );
  hadd1 \G1/G1_1(12)/U1_1 (
      .A(A[12]), .B(carry[12]), .S(SUM[12]), .CO(carry[13])
  );
  hadd1 \G1/G1_1(11)/U1_1 (
      .A(A[11]), .B(carry[11]), .S(SUM[11]), .CO(carry[12])
  );
  hadd1 \G1/G1_1(10)/U1_1 (
      .A(A[10]), .B(carry[10]), .S(SUM[10]), .CO(carry[11])
  );
  hadd1 \G1/G1_1(9)/U1_1 (
      .A(A[9]), .B(carry[9]), .S(SUM[9]), .CO(carry[10])
  );
  hadd1 \G1/G1_1(8)/U1_1 (
      .A(A[8]), .B(carry[8]), .S(SUM[8]), .CO(carry[9])
  );
  hadd1 \G1/G1_1(7)/U1_1 (
      .A(A[7]), .B(carry[7]), .S(SUM[7]), .CO(carry[8])
  );
  hadd1 \G1/G1_1(6)/U1_1 (
      .A(A[6]), .B(carry[6]), .S(SUM[6]), .CO(carry[7])
  );
  hadd1 \G1/G1_1(5)/U1_1 (
      .A(A[5]), .B(carry[5]), .S(SUM[5]), .CO(carry[6])
  );
  hadd1 \G1/G1_1(4)/U1_1 (
      .A(A[4]), .B(carry[4]), .S(SUM[4]), .CO(carry[5])
  );
  hadd1 \G1/G1_1(3)/U1_1 (
      .A(A[3]), .B(carry[3]), .S(SUM[3]), .CO(carry[4])
  );
  hadd1 \G1/G1_1(2)/U1_1 (
      .A(A[2]), .B(carry[2]), .S(SUM[2]), .CO(carry[3])
  );
  hadd1 \G1/G1_1(1)/U1_1 (
      .A(A[1]), .B(A[0]), .S(SUM[1]), .CO(carry[2])
  );
  inv02 U1(
      .A(A[0]), .Y(SUM[0])
  );
  xor02 U2(
      .A0(carry[31]), .A1(A[31]), .Y(SUM[31])
  );
endmodule

module clock_divider2(clk_i, rst_i, clk_o);
  input  clk_i, rst_i;
  output clk_o;

  wire [31:0] counter;
  wire N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
       N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
       N34, N35, N36, N37, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
       N54, N55, N61, N62, N63, N66, N67, N68, n15, n64, n1, n2, n3, n4, n5,
       n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17, n18, n19, n20, n21,
       n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
       n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
       n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
       n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
       n79, n80, n81, n82, n83, n84, n85, n86, n87, n88;

  dffr \counter_reg[0] (
      .D(N37), .CLK(clk_i), .R(n2), .Q(counter[0]), .QB()
  );
  dffr \counter_reg[1] (
      .D(n88), .CLK(clk_i), .R(n3), .Q(counter[1]), .QB()
  );
  dffr \counter_reg[2] (
      .D(n87), .CLK(clk_i), .R(n4), .Q(counter[2]), .QB()
  );
  dffr \counter_reg[3] (
      .D(n86), .CLK(clk_i), .R(n2), .Q(counter[3]), .QB()
  );
  dffr \counter_reg[4] (
      .D(n85), .CLK(clk_i), .R(n3), .Q(counter[4]), .QB()
  );
  dffr \counter_reg[5] (
      .D(n84), .CLK(clk_i), .R(n4), .Q(counter[5]), .QB()
  );
  dffr \counter_reg[6] (
      .D(n83), .CLK(clk_i), .R(n2), .Q(counter[6]), .QB()
  );
  dffr \counter_reg[7] (
      .D(N44), .CLK(clk_i), .R(n4), .Q(counter[7]), .QB()
  );
  dffr \counter_reg[8] (
      .D(N45), .CLK(clk_i), .R(n3), .Q(counter[8]), .QB()
  );
  dffr \counter_reg[9] (
      .D(N46), .CLK(clk_i), .R(n2), .Q(counter[9]), .QB()
  );
  dffr \counter_reg[10] (
      .D(N47), .CLK(clk_i), .R(n4), .Q(counter[10]), .QB(n15)
  );
  dffr \counter_reg[11] (
      .D(N48), .CLK(clk_i), .R(n3), .Q(counter[11]), .QB()
  );
  dffr \counter_reg[12] (
      .D(N49), .CLK(clk_i), .R(n2), .Q(counter[12]), .QB(n74)
  );
  dffr \counter_reg[13] (
      .D(N50), .CLK(clk_i), .R(n4), .Q(counter[13]), .QB(n75)
  );
  dffr \counter_reg[14] (
      .D(N51), .CLK(clk_i), .R(n3), .Q(counter[14]), .QB()
  );
  dffr \counter_reg[15] (
      .D(N52), .CLK(clk_i), .R(n2), .Q(counter[15]), .QB(n70)
  );
  dffr \counter_reg[16] (
      .D(N53), .CLK(clk_i), .R(n4), .Q(counter[16]), .QB(n71)
  );
  dffr \counter_reg[17] (
      .D(N54), .CLK(clk_i), .R(n3), .Q(counter[17]), .QB(n72)
  );
  dffr \counter_reg[18] (
      .D(N55), .CLK(clk_i), .R(n2), .Q(counter[18]), .QB()
  );
  dffr \counter_reg[19] (
      .D(n82), .CLK(clk_i), .R(n4), .Q(counter[19]), .QB()
  );
dffr \counter_reg[20] (
      .D(n81), .CLK(clk_i), .R(n3), .Q(counter[20]), .QB(n73)
  );
  dffr \counter_reg[21] (
      .D(n80), .CLK(clk_i), .R(n2), .Q(counter[21]), .QB(n66)
  );
  dffr \counter_reg[22] (
      .D(n79), .CLK(clk_i), .R(n3), .Q(counter[22]), .QB()
  );
  dffr \counter_reg[23] (
      .D(n78), .CLK(clk_i), .R(n4), .Q(counter[23]), .QB(n67)
  );
  dffr \counter_reg[24] (
      .D(N61), .CLK(clk_i), .R(n1), .Q(counter[24]), .QB(n68)
  );
  dffr \counter_reg[25] (
      .D(N62), .CLK(clk_i), .R(n1), .Q(counter[25]), .QB(n69)
  );
  dffr \counter_reg[26] (
      .D(N63), .CLK(clk_i), .R(n1), .Q(counter[26]), .QB()
  );
  dffr \counter_reg[27] (
      .D(n77), .CLK(clk_i), .R(n1), .Q(counter[27]), .QB()
  );
  dffr \counter_reg[28] (
      .D(n76), .CLK(clk_i), .R(n1), .Q(counter[28]), .QB()
  );
  dffr \counter_reg[29] (
      .D(N66), .CLK(clk_i), .R(n1), .Q(counter[29]), .QB()
  );
  dffr \counter_reg[30] (
      .D(N67), .CLK(clk_i), .R(n1), .Q(counter[30]), .QB()
  );
  dffr \counter_reg[31] (
      .D(N68), .CLK(clk_i), .R(n1), .Q(counter[31]), .QB()
  );
  dffr clk_o_reg(
      .D(n64), .CLK(clk_i), .R(n1), .Q(clk_o), .QB()
  );
  clock_divider_DW01_inc_0 add_42(
      .A(counter), .SUM({N36, N35, N34, N33, N32, N31, N30, N29, N28, N27,
      N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13,
      N12, N11, N10, N9, N8, N7, N6, N5})
  );
  inv02 U3(
      .A(rst_i), .Y(n1)
  );
  inv01 U4(
      .A(rst_i), .Y(n2)
  );
  inv01 U5(
      .A(rst_i), .Y(n3)
  );
  inv01 U6(
      .A(rst_i), .Y(n4)
  );
  and04 U7(
      .A0(n55), .A1(n56), .A2(n57), .A3(n58), .Y(n45)
  );
  inv02 U8(
      .A(n45), .Y(n5)
  );
  inv01 U9(
      .A(n45), .Y(n6)
  );
  inv01 U10(
      .A(n45), .Y(n7)
  );
  inv01 U11(
      .A(n45), .Y(n8)
  );
  inv01 U12(
      .A(n9), .Y(n79)
  );
  inv01 U13(
      .A(n10), .Y(n80)
  );
  inv01 U14(
      .A(n11), .Y(n81)
  );
  inv01 U15(
      .A(n12), .Y(n82)
  );
  mux21 U16(
      .A0(n13), .A1(clk_o), .S0(n14), .Y(n64)
  );
  nor02ii U17(
      .A0(n16), .A1(n13), .Y(n14)
  );
  nor04 U18(
      .A0(n17), .A1(n18), .A2(n19), .A3(n20), .Y(n16)
  );
  nand04 U19(
      .A0(N13), .A1(N15), .A2(N12), .A3(n21), .Y(n20)
  );
  nor02 U20(
      .A0(n22), .A1(n10), .Y(n21)
  );
  nand04 U21(
      .A0(n23), .A1(n24), .A2(N10), .A3(n25), .Y(n19)
  );
  nor03 U22(
      .A0(n26), .A1(n27), .A2(n28), .Y(n25)
  );
  inv01 U23(
      .A(N14), .Y(n24)
  );
  or04 U24(
      .A0(N17), .A1(N19), .A2(N16), .A3(n29), .Y(n18)
  );
  or03 U25(
      .A0(N20), .A1(N24), .A2(N21), .Y(n29)
  );
  nand04 U26(
      .A0(n30), .A1(n31), .A2(n32), .A3(n33), .Y(n17)
  );
  nor03 U27(
      .A0(N7), .A1(N9), .A2(N8), .Y(n33)
  );
 inv01 U28(
      .A(N25), .Y(n32)
  );
  nand04 U29(
      .A0(n34), .A1(n35), .A2(n36), .A3(n37), .Y(n13)
  );
  nor04 U30(
      .A0(n38), .A1(n39), .A2(N37), .A3(n22), .Y(n37)
  );
  nand04 U31(
      .A0(n40), .A1(n41), .A2(n42), .A3(n43), .Y(n22)
  );
  nor04 U32(
      .A0(n44), .A1(n78), .A2(n76), .A3(n77), .Y(n43)
  );
  and02 U33(
      .A0(N32), .A1(n5), .Y(n77)
  );
  and02 U34(
      .A0(N33), .A1(n5), .Y(n76)
  );
  and02 U35(
      .A0(N28), .A1(n7), .Y(n78)
  );
  nand02 U36(
      .A0(n46), .A1(n9), .Y(n44)
  );
  nand02 U37(
      .A0(N27), .A1(n6), .Y(n9)
  );
  nor03 U38(
      .A0(N63), .A1(N67), .A2(N66), .Y(n42)
  );
  nand03 U39(
      .A0(n47), .A1(n48), .A2(n49), .Y(n39)
  );
  nand04 U40(
      .A0(n50), .A1(n51), .A2(n52), .A3(n53), .Y(n38)
  );
  nor03 U41(
      .A0(N50), .A1(N52), .A2(N51), .Y(n53)
  );
  nor04 U42(
      .A0(n54), .A1(n85), .A2(n83), .A3(n84), .Y(n36)
  );
  and02 U43(
      .A0(N10), .A1(n8), .Y(n84)
  );
  nor02ii U44(
      .A0(n23), .A1(n8), .Y(n83)
  );
  inv01 U45(
      .A(N11), .Y(n23)
  );
  and02 U46(
      .A0(N9), .A1(n6), .Y(n85)
  );
  nand03 U47(
      .A0(n11), .A1(n10), .A2(n12), .Y(n54)
  );
 nand02 U48(
      .A0(N24), .A1(n7), .Y(n12)
  );
  nand02 U49(
      .A0(N26), .A1(n8), .Y(n10)
  );
  nand02 U50(
      .A0(N25), .A1(n6), .Y(n11)
  );
  nor03 U51(
      .A0(n88), .A1(n86), .A2(n87), .Y(n35)
  );
  and02 U52(
      .A0(N7), .A1(n7), .Y(n87)
  );
  and02 U53(
      .A0(N8), .A1(n5), .Y(n86)
  );
  nor02ii U54(
      .A0(n31), .A1(n6), .Y(n88)
  );
  inv01 U55(
      .A(N6), .Y(n31)
  );
  nor03 U56(
      .A0(N53), .A1(N55), .A2(N54), .Y(n34)
  );
  inv01 U57(
      .A(n46), .Y(N68)
  );
  nand02 U58(
      .A0(N36), .A1(n7), .Y(n46)
  );
  and02 U59(
      .A0(N35), .A1(n5), .Y(N67)
  );
  and02 U60(
      .A0(N34), .A1(n5), .Y(N66)
  );
  and02 U61(
      .A0(N31), .A1(n5), .Y(N63)
  );
  inv01 U62(
      .A(n41), .Y(N62)
  );
  nand02 U63(
      .A0(N30), .A1(n8), .Y(n41)
  );
  inv01 U64(
      .A(n40), .Y(N61)
  );
  nand02 U65(
      .A0(N29), .A1(n6), .Y(n40)
  );
  nor02ii U66(
      .A0(n27), .A1(n7), .Y(N55)
  );
  inv01 U67(
      .A(N23), .Y(n27)
  );
 nor02ii U68(
      .A0(n28), .A1(n8), .Y(N54)
  );
  inv01 U69(
      .A(N22), .Y(n28)
  );
  and02 U70(
      .A0(N21), .A1(n5), .Y(N53)
  );
  and02 U71(
      .A0(N20), .A1(n5), .Y(N52)
  );
  and02 U72(
      .A0(n8), .A1(N19), .Y(N51)
  );
  nor02ii U73(
      .A0(n26), .A1(n6), .Y(N50)
  );
  inv01 U74(
      .A(N18), .Y(n26)
  );
  inv01 U75(
      .A(n51), .Y(N49)
  );
  nand02 U76(
      .A0(N17), .A1(n7), .Y(n51)
  );
  inv01 U77(
      .A(n50), .Y(N48)
  );
  nand02 U78(
      .A0(N16), .A1(n8), .Y(n50)
  );
  inv01 U79(
      .A(n52), .Y(N47)
  );
  nand02 U80(
      .A0(N15), .A1(n6), .Y(n52)
  );
  inv01 U81(
      .A(n48), .Y(N46)
  );
  nand02 U82(
      .A0(N14), .A1(n7), .Y(n48)
  );
  inv01 U83(
      .A(n47), .Y(N45)
  );
  nand02 U84(
      .A0(N13), .A1(n8), .Y(n47)
  );
  inv01 U85(
      .A(n49), .Y(N44)
  );
  nand02 U86(
      .A0(N12), .A1(n6), .Y(n49)
  );
  nor02ii U87(
      .A0(n30), .A1(n7), .Y(N37)
  );
 inv01 U88(
      .A(N5), .Y(n30)
  );
  nor04 U89(
      .A0(n59), .A1(n60), .A2(n61), .A3(n62), .Y(n58)
  );
  nand04 U90(
      .A0(n74), .A1(n75), .A2(n15), .A3(counter[3]), .Y(n62)
  );
  nand04 U91(
      .A0(counter[2]), .A1(counter[22]), .A2(counter[1]), .A3(counter[9]), .Y(n61)
  );
  nand04 U92(
      .A0(counter[8]), .A1(counter[5]), .A2(counter[4]), .A3(counter[0]), .Y(n60)
  );
  nand04 U93(
      .A0(counter[19]), .A1(counter[18]), .A2(counter[14]), .A3(counter[11]), .Y(n59)
  );
  nor02 U94(
      .A0(n63), .A1(n65), .Y(n57)
  );
  nand04 U95(
      .A0(n66), .A1(n67), .A2(n68), .A3(n69), .Y(n65)
  );
  nand04 U96(
      .A0(n70), .A1(n71), .A2(n72), .A3(n73), .Y(n63)
  );
  nor04 U97(
      .A0(counter[29]), .A1(counter[28]), .A2(counter[27]), .A3(counter[26]), .Y(n56)
  );
  nor04 U98(
      .A0(counter[7]), .A1(counter[6]), .A2(counter[31]), .A3(counter[30]), .Y(n55)
  );
endmodule

